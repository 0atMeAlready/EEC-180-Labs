module RAM (

    input [3:0] Address, Data_in,
    input Write_Enable, Clock,
    output [3:0] Data_out

)

reg [3:0] memory [15:0] /*synthesis ramstyle = "M9K" */

always @ (posedge clk) begin

    if (mwr) 
    
    memory [addr] <= mdi; //writes memory
    mdo <= memory [addr]; //reads memory

end

endmodule

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module partI(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,
	output		     [7:0]		HEX2,
	output		     [7:0]		HEX3,
	output		     [7:0]		HEX4,
	output		     [7:0]		HEX5,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================
wire Enable, RAM_SELECT, CLK, Add, Data_in, RAM1_OUT, RAM0_OUT;

//=======================================================
//  Structural coding
//=======================================================
assign Enable = SW[9];
assign RAM_SELECT = SW[8];
assign CLK = KEY[0];
assign Add = SW[7:4];
assign Data_in = SW[3:0];

// Generate write enable signals for RAM0 and RAM1
wire RAM0_WE = Write_Enable & ~RAM_SELECT;  // Write to RAM0 when RAM_SELECT = 0
wire RAM1_WE = Write_Enable &  RAM_SELECT;  // Write to RAM1 when RAM_SELECT = 1

// Instantiate RAM0
RAM RAM0 (
    .Address(Address),
    .Data_in(Data_in),
    .Write_Enable(RAM0_WE),
    .Clock(CLK),
    .Data_out(RAM0_OUT)
);

// Instantiate RAM1
RAM RAM1 (
    .Address(Address),
    .Data_in(Data_in),
    .Write_Enable(RAM1_WE),
    .Clock(CLK),
    .Data_out(RAM1_OUT)
);

//=======================================================
//  Display Output Mapping
//=======================================================

// Display Address on HEX3
hex_decoder hex3_inst (
    .binary_in(Address),
    .seg_out(HEX3)
);

// Display Data_in on HEX2
hex_decoder hex2_inst (
    .binary_in(Data_in),
    .seg_out(HEX2)
);

// Display RAM1 output on HEX1
hex_decoder hex1_inst (
    .binary_in(RAM1_OUT),
    .seg_out(HEX1)
);

// Display RAM0 output on HEX0
hex_decoder hex0_inst (
    .binary_in(RAM0_OUT),
    .seg_out(HEX0)
);

endmodule