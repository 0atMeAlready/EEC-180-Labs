module RAM (
<<<<<<< HEAD

    input [3:0] Address, Data_in,
    input Write_Enable, Clock,
    output [3:0] Data_out

)

reg [3:0] memory [15:0] /*synthesis ramstyle = "M9K" */

always @ (posedge clk) begin

    if (mwr) 
    
    memory [addr] <= mdi; //writes memory
    mdo <= memory [addr]; //reads memory

end

endmodule

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module partI(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,
	output		     [7:0]		HEX2,
	output		     [7:0]		HEX3,
	output		     [7:0]		HEX4,
	output		     [7:0]		HEX5,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================
wire Enable, RAM_SELECT, CLK, Add, Data_in, RAM1_OUT, RAM0_OUT;

//=======================================================
//  Structural coding
//=======================================================
assign Enable = SW[9];
assign RAM_SELECT = SW[8];
assign CLK = KEY[0];
assign Add = SW[7:4];
assign Data_in = SW[3:0];

// Generate write enable signals for RAM0 and RAM1
wire RAM0_WE = Write_Enable & ~RAM_SELECT;  // Write to RAM0 when RAM_SELECT = 0
wire RAM1_WE = Write_Enable &  RAM_SELECT;  // Write to RAM1 when RAM_SELECT = 1

// Instantiate RAM0
RAM RAM0 (
    .Address(Address),
    .Data_in(Data_in),
    .Write_Enable(RAM0_WE),
    .Clock(CLK),
    .Data_out(RAM0_OUT)
);

// Instantiate RAM1
RAM RAM1 (
    .Address(Address),
    .Data_in(Data_in),
    .Write_Enable(RAM1_WE),
    .Clock(CLK),
    .Data_out(RAM1_OUT)
);

//=======================================================
//  Display Output Mapping
//=======================================================

// Display Address on HEX3
hex_decoder hex3_inst (
    .binary_in(Address),
    .seg_out(HEX3)
);

// Display Data_in on HEX2
hex_decoder hex2_inst (
    .binary_in(Data_in),
    .seg_out(HEX2)
);

// Display RAM1 output on HEX1
hex_decoder hex1_inst (
    .binary_in(RAM1_OUT),
    .seg_out(HEX1)
);

// Display RAM0 output on HEX0
hex_decoder hex0_inst (
    .binary_in(RAM0_OUT),
    .seg_out(HEX0)
);

endmodule
=======
    input wire [3:0] Addr,
    input wire [7:0] MDI,
    input wire Write_Enable, CLK,
    output reg [7:0] MDO
);
    reg [7:0] memory [15:0];
    always @(posedge CLK) begin
        if (Write_Enable)
            memory[Addr] <= MDI;
        MDO <= memory[Addr];
    end
endmodule

module SquareRoot (
    input wire CLK, ResetN, St,
    input wire [7:0] N,
    output reg Done,
    output reg [3:0] Sqrt
);
    reg [7:0] R;
    reg [3:0] count;
    reg [7:0] odd;
    reg calculating;
    
    always @(posedge CLK or negedge ResetN) begin
        if (!ResetN) begin
            Sqrt <= 4'b0;
            Done <= 0;
            calculating <= 0;
        end 
        else if (St && !calculating) begin
            R <= N;
            odd <= 8'd1;
            count <= 4'b0;
            Done <= 0;
            calculating <= 1;
        end 
        else if (calculating) begin
            if (R >= odd) begin
                R <= R - odd;
                odd <= odd + 8'd2;
                count <= count + 1;
            end else begin
                Sqrt <= count;
                Done <= 1;
                calculating <= 0;
            end
        end
    end
endmodule

module Controller (
    input wire CLK, ResetN, St,
    output wire Done,
    output wire [3:0] Sqrt,
    output wire [7:0] N
);
    reg [3:0] Addr;
    reg Write_Enable;
    wire [7:0] MDO;
    wire [3:0] Sqrt_Result;
    reg Output_Write_Enable;
    reg [3:0] Out_Addr;
    
    RAM ram_inst (
        .Addr(Addr),
        .MDI(8'b0),
        .Write_Enable(Write_Enable),
        .CLK(CLK),
        .MDO(MDO)
    );
    
    SquareRoot sqrt_inst (
        .CLK(CLK),
        .ResetN(ResetN),
        .St(St),
        .N(MDO),
        .Done(Done),
        .Sqrt(Sqrt_Result)
    );
    
    RAM output_ram (
        .Addr(Out_Addr),
        .MDI({4'b0, Sqrt_Result}),
        .Write_Enable(Output_Write_Enable),
        .CLK(CLK),
        .MDO()
    );
    
    assign N = MDO;
    assign Sqrt = Sqrt_Result;
    
    always @(posedge CLK or negedge ResetN) begin
        if (!ResetN) begin
            Addr <= 0;
            Write_Enable <= 1;
            Out_Addr <= 0;
            Output_Write_Enable <= 0;
        end 
        else if (St) begin
            if (Addr == 4'b1111) begin
                Addr <= 0;
                Write_Enable <= 0;
            end else begin
                Addr <= Addr + 1;
            end
            if (Done) begin
                Output_Write_Enable <= 1;
                Out_Addr <= Addr;
            end else begin
                Output_Write_Enable <= 0;
            end
        end
    end
endmodule

module tb_sqrt;
    parameter num_vectors = 16;
    reg CLK, ResetN, St;
    wire Done;
    reg [7:0] MDI;
    wire [3:0] Sqrt;
    reg [7:0] vectors [0:num_vectors-1];
    integer i;
    wire [7:0] MDO_wire;
    reg [3:0] Addr;
    reg Write_Enable;
    
    RAM ram_inst (
        .Addr(Addr),
        .MDI(MDI),
        .Write_Enable(Write_Enable),
        .CLK(CLK),
        .MDO(MDO_wire)
    );
    
    SquareRoot sqrt_inst (
        .CLK(CLK),
        .ResetN(ResetN),
        .St(St),
        .N(MDO_wire),
        .Done(Done),
        .Sqrt(Sqrt)
    );
    
    Controller UUT (
        .CLK(CLK),
        .ResetN(ResetN),
        .St(St),
        .Done(Done),
        .Sqrt(Sqrt),
        .N(MDO_wire)
    );
    
    initial begin
        CLK = 0;
        forever #20 CLK = ~CLK;
    end
    
    initial begin
        ResetN = 0;
        St = 0;
        #80 ResetN = 1;
        $readmemb("testvecs", vectors);
        for (i = 0; i < num_vectors; i = i + 1) begin
            MDI = vectors[i];
            #20 St = 1;
            wait (Done == 1);
            $display("Input=0x%h, SqRt=0x%h", MDI, Sqrt);
            #20 St = 0;
            wait (Done == 0);
        end
        $finish;
    end
endmodule
>>>>>>> e459053b692d03062a2895e52efafc5c956584d3
